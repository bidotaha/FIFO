package shared_pkg ;

bit test_finished ;

int error_count = 0 ;
int correct_count = 0 ;
endpackage